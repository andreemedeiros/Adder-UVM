interface fulladder_if(input sig_clk,sig_rst);
  logic sig_a;
  logic sig_b;
  logic sig_c_in;
  logic sig_sum;
  logic sig_c_out;
endinterface