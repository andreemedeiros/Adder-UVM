package full_add_pkg;
import uvm_pkg::*;
`include "full_adder_seq_item.sv"
`include "full_add_sequencer.sv"
`include "full_add_driver.sv"
`include "full_add_monitor.sv"
`include "full_adder_agent.sv"
`include "full_add_env.sv"
`include "full_adder_seq.sv"
`include "full_add_test.sv"
endpackage