package pkg;
import uvm_pkg::*;
`include "adder_seq_item.sv"
`include "add_sequencer.sv"
`include "add_driver.sv"
`include "add_monitor.sv"
`include "adder_agent.sv"
`include "add_env.sv"
`include "adder_seq.sv"
`include "add_test.sv"
endpackage
