package full_add_pkg;
import uvm_pkg::*;
`include "seq_item.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "env.sv"
`include "seq.sv"
`include "test.sv"
endpackage